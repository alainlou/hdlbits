module top_module ( input a, input b, output out );
    mod_a block ( a, b, out );
endmodule
